// Uncomment to flip on the debug ILAs
//`define USING_DEBUG 1