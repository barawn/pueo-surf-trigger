package pueo_beams;
	localparam TRIPLET_ADDER_TOTAL = 67;
	localparam DOUBLET_ADDER_TOTAL = 12;
	localparam NUM_BEAMS = 46;

	localparam int TRIPLET_ADDER_INDICES [0:TRIPLET_ADDER_TOTAL-1][0:2] = '{
		'{ 1,3,5 } ,
		'{ 5,6,7 } ,
		'{ 1,6,7 } ,
		'{ 1,5,6 } ,
		'{ 1,2,3 } ,
		'{ 1,3,6 } ,
		'{ 1,2,3 } ,
		'{ 3,5,7 } ,
		'{ 2,3,5 } ,
		'{ 2,3,7 } ,
		'{ 1,2,7 } ,
		'{ 2,6,7 } ,
		'{ 2,5,7 } ,
		'{ 1,3,6 } ,
		'{ 5,6,7 } ,
		'{ 5,6,7 } ,
		'{ 1,6,7 } ,
		'{ 3,5,6 } ,
		'{ 2,3,6 } ,
		'{ 2,3,5 } ,
		'{ 1,2,3 } ,
		'{ 2,5,7 } ,
		'{ 5,6,7 } ,
		'{ 1,3,6 } ,
		'{ 1,2,3 } ,
		'{ 1,3,6 } ,
		'{ 1,2,3 } ,
		'{ 1,6,7 } ,
		'{ 1,2,7 } ,
		'{ 3,5,6 } ,
		'{ 1,2,6 } ,
		'{ 1,2,3 } ,
		'{ 1,2,6 } ,
		'{ 5,6,7 } ,
		'{ 1,2,7 } ,
		'{ 3,5,6 } ,
		'{ 1,5,7 } ,
		'{ 5,6,7 } ,
		'{ 1,2,7 } ,
		'{ 5,6,7 } ,
		'{ 2,5,7 } ,
		'{ 2,5,7 } ,
		'{ 1,2,3 } ,
		'{ 5,6,7 } ,
		'{ 1,2,3 } ,
		'{ 5,6,7 } ,
		'{ 1,2,5 } ,
		'{ 1,2,3 } ,
		'{ 3,6,7 } ,
		'{ 5,6,7 } ,
		'{ 5,6,7 } ,
		'{ 3,5,6 } ,
		'{ 1,2,3 } ,
		'{ 1,5,7 } ,
		'{ 1,2,3 } ,
		'{ 3,5,7 } ,
		'{ 1,2,3 } ,
		'{ 2,3,6 } ,
		'{ 2,5,7 } ,
		'{ 5,6,7 } ,
		'{ 1,2,3 } ,
		'{ 3,5,7 } ,
		'{ 2,6,7 } ,
		'{ 5,6,7 } ,
		'{ 5,6,7 } ,
		'{ 1,2,3 } ,
		'{ 1,2,3 }  };

	localparam int TRIPLET_ADDER_DELAYS [0:TRIPLET_ADDER_TOTAL-1][0:2] = '{
		'{ 30,38,30 } ,
		'{ 10,10,9 } ,
		'{ 28,31,35 } ,
		'{ 29,28,32 } ,
		'{ 4,2,0 } ,
		'{ 11,10,10 } ,
		'{ 11,11,11 } ,
		'{ 42,32,42 } ,
		'{ 31,35,28 } ,
		'{ 33,37,36 } ,
		'{ 21,23,27 } ,
		'{ 34,34,38 } ,
		'{ 39,34,44 } ,
		'{ 6,3,5 } ,
		'{ 21,23,25 } ,
		'{ 12,12,12 } ,
		'{ 27,32,36 } ,
		'{ 15,13,14 } ,
		'{ 37,41,36 } ,
		'{ 16,17,17 } ,
		'{ 25,29,32 } ,
		'{ 4,7,4 } ,
		'{ 26,30,33 } ,
		'{ 7,4,4 } ,
		'{ 13,13,13 } ,
		'{ 34,44,39 } ,
		'{ 25,28,31 } ,
		'{ 16,18,18 } ,
		'{ 22,24,26 } ,
		'{ 26,22,24 } ,
		'{ 23,25,25 } ,
		'{ 8,7,6 } ,
		'{ 32,37,37 } ,
		'{ 25,28,31 } ,
		'{ 15,15,14 } ,
		'{ 27,21,23 } ,
		'{ 16,15,16 } ,
		'{ 17,18,19 } ,
		'{ 13,14,15 } ,
		'{ 9,8,7 } ,
		'{ 5,6,3 } ,
		'{ 10,11,10 } ,
		'{ 27,31,34 } ,
		'{ 5,3,1 } ,
		'{ 9,9,8 } ,
		'{ 8,7,6 } ,
		'{ 15,16,15 } ,
		'{ 17,18,19 } ,
		'{ 16,16,16 } ,
		'{ 19,21,23 } ,
		'{ 18,19,20 } ,
		'{ 14,15,15 } ,
		'{ 9,8,7 } ,
		'{ 32,32,40 } ,
		'{ 20,22,24 } ,
		'{ 28,23,28 } ,
		'{ 18,19,20 } ,
		'{ 17,17,15 } ,
		'{ 11,10,9 } ,
		'{ 13,13,13 } ,
		'{ 5,3,1 } ,
		'{ 41,32,41 } ,
		'{ 34,35,39 } ,
		'{ 4,2,0 } ,
		'{ 24,27,30 } ,
		'{ 23,26,29 } ,
		'{ 19,21,23 }  };

	localparam int DOUBLET_ADDER_INDICES [0:DOUBLET_ADDER_TOTAL-1][0:1] = '{
		'{ 0,4  } ,
		'{ 0,4  } ,
		'{ 0,4  } ,
		'{ 0,4  } ,
		'{ 0,4  } ,
		'{ 0,4  } ,
		'{ 0,4  } ,
		'{ 0,4  } ,
		'{ 0,4  } ,
		'{ 0,4  } ,
		'{ 0,4  } ,
		'{ 0,4  }  };

	localparam int DOUBLET_ADDER_DELAYS [0:DOUBLET_ADDER_TOTAL-1][0:1] = '{
		'{ 1,1  } ,
		'{ 1,2  } ,
		'{ 3,0  } ,
		'{ 1,0  } ,
		'{ 1,4  } ,
		'{ 2,0  } ,
		'{ 4,0  } ,
		'{ 0,1  } ,
		'{ 0,3  } ,
		'{ 5,1  } ,
		'{ 0,2  } ,
		'{ 0,0  }  };

	localparam int BEAM_CONTENTS [0:NUM_BEAMS-1][0:2] = '{
		'{ 4,63,4 } ,
		'{ 40,13,4 } ,
		'{ 31,45,4 } ,
		'{ 52,39,7 } ,
		'{ 41,5,7 } ,
		'{ 24,59,7 } ,
		'{ 48,46,0 } ,
		'{ 37,47,0 } ,
		'{ 66,49,0 } ,
		'{ 28,29,0 } ,
		'{ 55,30,3 } ,
		'{ 33,26,3 } ,
		'{ 2,8,2 } ,
		'{ 11,0,2 } ,
		'{ 61,32,6 } ,
		'{ 12,25,6 } ,
		'{ 4,43,8 } ,
		'{ 13,21,8 } ,
		'{ 39,31,8 } ,
		'{ 44,1,10 } ,
		'{ 6,15,10 } ,
		'{ 38,51,10 } ,
		'{ 19,27,0 } ,
		'{ 50,47,11 } ,
		'{ 14,54,0 } ,
		'{ 10,29,3 } ,
		'{ 65,64,3 } ,
		'{ 20,22,3 } ,
		'{ 16,8,5 } ,
		'{ 0,62,5 } ,
		'{ 7,32,2 } ,
		'{ 60,63,8 } ,
		'{ 23,40,1 } ,
		'{ 52,45,1 } ,
		'{ 5,58,1 } ,
		'{ 24,15,1 } ,
		'{ 17,34,0 } ,
		'{ 57,36,11 } ,
		'{ 37,56,11 } ,
		'{ 54,49,3 } ,
		'{ 28,35,3 } ,
		'{ 64,26,5 } ,
		'{ 42,22,2 } ,
		'{ 3,9,2 } ,
		'{ 53,18,9 } ,
		'{ 12,25,9 }  };

	localparam TRIPLET_DUMMY_TOTAL = 4;
	localparam DOUBLET_DUMMY_TOTAL = 2;
	localparam NUM_BEAMS_DUMMY = 2;

	localparam int TRIPLET_DUMMY_DELAYS [0:TRIPLET_DUMMY_TOTAL-1][0:2] = '{
		'{0,0,0},
		'{0,0,0},
		'{11,11,11},
		'{12,12,12} };

	localparam int TRIPLET_DUMMY_INDICES [0:TRIPLET_DUMMY_TOTAL-1][0:2] = '{
		'{1,2,3},
		'{5,6,7},
		'{1,2,3},
		'{5,6,7} };

	localparam int DOUBLET_DUMMY_DELAYS [0:DOUBLET_DUMMY_TOTAL-1][0:1] = '{
		'{0,0},
		'{0,2} };

	localparam int BEAM_CONTENTS_DUMMY [0:NUM_BEAMS_DUMMY-1] = '{
		'{0,1,0},
		'{2,3,1} };

endpackage
