// Uncomment to use the debug pathways in the trigger
//`define USING_DEBUG 0