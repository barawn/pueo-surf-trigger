`ifndef PUEO_BEAMS_SV
`define PUEO_BEAMS_SV

// Vivado won't show 
package pueo_beams;
	localparam int NUM_BEAM = 48;

	localparam int SAMPLE_STORE_DEPTH = 4;

	localparam int LEFT_ADDER_LEN = 7;

	localparam int LEFT_STORE_DEPTH = 2;

	localparam int RIGHT_ADDER_LEN = 7;

	localparam int RIGHT_STORE_DEPTH = 2;

	localparam int TOP_ADDER_LEN = 5;

	localparam int TOP_STORE_DEPTH = 1;

	localparam int META0_INDICES [0:21] = '{
		18,
		19,
		20,
		25,
		26,
		27,
		32,
		33,
		34,
		46,
		47,
		255,
		255,
		255,
		255,
		255,
		255,
		255,
		255,
		255,
		255,
		255 };


	localparam int META1_INDICES [0:21] = '{
		4,
		5,
		6,
		11,
		12,
		13,
		18,
		19,
		20,
		39,
		40,
		41,
		255,
		255,
		255,
		255,
		255,
		255,
		255,
		255,
		255,
		255 };


	localparam int META2_INDICES [0:21] = '{
		17,
		18,
		19,
		24,
		25,
		26,
		31,
		32,
		33,
		45,
		46,
		47,
		255,
		255,
		255,
		255,
		255,
		255,
		255,
		255,
		255,
		255 };


	localparam int META3_INDICES [0:21] = '{
		3,
		4,
		5,
		10,
		11,
		12,
		17,
		18,
		19,
		38,
		39,
		40,
		255,
		255,
		255,
		255,
		255,
		255,
		255,
		255,
		255,
		255 };


	localparam int META4_INDICES [0:21] = '{
		15,
		16,
		17,
		22,
		23,
		24,
		29,
		30,
		31,
		43,
		44,
		45,
		255,
		255,
		255,
		255,
		255,
		255,
		255,
		255,
		255,
		255 };


	localparam int META5_INDICES [0:21] = '{
		1,
		2,
		3,
		8,
		9,
		10,
		15,
		16,
		17,
		36,
		37,
		38,
		255,
		255,
		255,
		255,
		255,
		255,
		255,
		255,
		255,
		255 };


	localparam int META6_INDICES [0:21] = '{
		14,
		15,
		16,
		21,
		22,
		23,
		28,
		29,
		30,
		42,
		43,
		44,
		255,
		255,
		255,
		255,
		255,
		255,
		255,
		255,
		255,
		255 };


	localparam int META7_INDICES [0:21] = '{
		0,
		1,
		2,
		7,
		8,
		9,
		14,
		15,
		16,
		35,
		36,
		37,
		255,
		255,
		255,
		255,
		255,
		255,
		255,
		255,
		255,
		255 };


	localparam int LEFT_ADDERS [0:6][0:2] = '{
		'{ 19,21,23 },
		'{ 9,9,9 },
		'{ 17,18,20 },
		'{ 1,0,0 },
		'{ 0,2,5 },
		'{ 13,14,15 },
		'{ 11,11,12 } };


	localparam int RIGHT_ADDERS [0:6][0:2] = '{
		'{ 16,18,20 },
		'{ 10,10,10 },
		'{ 15,16,18 },
		'{ 1,0,0 },
		'{ 0,2,5 },
		'{ 14,15,16 },
		'{ 12,12,13 } };


	localparam int TOP_ADDERS [0:4][0:1] = '{
		'{ 0,1 },
		'{ 0,0 },
		'{ 2,0 },
		'{ 0,2 },
		'{ 1,0 } };


	localparam int BEAM_INDICES [0:47][0:2] = '{
		'{ 1,1,3 },
		'{ 1,1,3 },
		'{ 1,1,0 },
		'{ 1,1,0 },
		'{ 1,1,0 },
		'{ 1,1,1 },
		'{ 1,1,1 },
		'{ 6,6,3 },
		'{ 6,6,3 },
		'{ 6,6,0 },
		'{ 6,6,1 },
		'{ 6,6,1 },
		'{ 6,6,4 },
		'{ 6,6,4 },
		'{ 5,5,3 },
		'{ 5,5,0 },
		'{ 5,5,0 },
		'{ 5,5,1 },
		'{ 5,5,1 },
		'{ 5,5,4 },
		'{ 5,5,4 },
		'{ 2,2,3 },
		'{ 2,2,0 },
		'{ 2,2,1 },
		'{ 2,2,1 },
		'{ 2,2,4 },
		'{ 2,2,4 },
		'{ 2,2,2 },
		'{ 0,0,0 },
		'{ 0,0,1 },
		'{ 0,0,1 },
		'{ 0,0,4 },
		'{ 0,0,4 },
		'{ 0,0,2 },
		'{ 0,0,2 },
		'{ 3,3,255 },
		'{ 3,3,255 },
		'{ 3,3,255 },
		'{ 3,3,255 },
		'{ 3,3,255 },
		'{ 3,3,255 },
		'{ 3,3,255 },
		'{ 4,4,255 },
		'{ 4,4,255 },
		'{ 4,4,255 },
		'{ 4,4,255 },
		'{ 4,4,255 },
		'{ 4,4,255 } };


	localparam int BEAM_LEFT_OFFSETS [0:47] = '{
		4,
		5,
		4,
		3,
		3,
		2,
		0,
		4,
		4,
		4,
		3,
		3,
		2,
		0,
		4,
		3,
		4,
		3,
		3,
		2,
		0,
		1,
		2,
		2,
		1,
		2,
		1,
		0,
		0,
		1,
		1,
		1,
		1,
		1,
		0,
		3,
		2,
		1,
		0,
		0,
		0,
		0,
		3,
		2,
		1,
		0,
		0,
		0 };


	localparam int BEAM_RIGHT_OFFSETS [0:47] = '{
		0,
		2,
		2,
		2,
		3,
		3,
		2,
		0,
		1,
		2,
		2,
		3,
		3,
		2,
		0,
		0,
		2,
		2,
		3,
		3,
		2,
		0,
		2,
		3,
		3,
		5,
		5,
		5,
		0,
		2,
		3,
		4,
		5,
		6,
		6,
		0,
		0,
		0,
		0,
		1,
		2,
		3,
		0,
		0,
		0,
		0,
		1,
		2 };


	localparam int BEAM_TOP_OFFSETS [0:47] = '{
		0,
		0,
		0,
		0,
		0,
		0,
		0,
		0,
		0,
		0,
		0,
		0,
		0,
		0,
		0,
		0,
		0,
		0,
		0,
		0,
		0,
		0,
		0,
		0,
		0,
		0,
		0,
		0,
		0,
		0,
		0,
		0,
		0,
		0,
		0,
		0,
		0,
		0,
		0,
		0,
		0,
		0,
		0,
		0,
		0,
		0,
		0,
		0 };


endpackage

`endif
