`define TRIPLET_ADDER_TOTAL 67
`define DOUBLET_ADDER_TOTAL 12
`define NUM_BEAM 46
`define TRIPLET_ADDER_INDICES '{ \
 '{ 2,5,7 } , \
 '{ 1,2,7 } , \
 '{ 1,5,7 } , \
 '{ 1,2,3 } , \
 '{ 5,6,7 } , \
 '{ 2,3,6 } , \
 '{ 1,2,3 } , \
 '{ 1,2,3 } , \
 '{ 1,2,5 } , \
 '{ 1,5,6 } , \
 '{ 1,2,3 } , \
 '{ 2,3,5 } , \
 '{ 3,5,6 } , \
 '{ 1,6,7 } , \
 '{ 1,5,7 } , \
 '{ 1,3,6 } , \
 '{ 1,2,6 } , \
 '{ 1,3,6 } , \
 '{ 1,2,3 } , \
 '{ 5,6,7 } , \
 '{ 1,2,3 } , \
 '{ 2,6,7 } , \
 '{ 5,6,7 } , \
 '{ 1,2,3 } , \
 '{ 5,6,7 } , \
 '{ 5,6,7 } , \
 '{ 1,2,3 } , \
 '{ 1,2,3 } , \
 '{ 1,2,6 } , \
 '{ 1,2,7 } , \
 '{ 2,5,7 } , \
 '{ 5,6,7 } , \
 '{ 1,6,7 } , \
 '{ 3,5,6 } , \
 '{ 2,5,7 } , \
 '{ 5,6,7 } , \
 '{ 1,3,5 } , \
 '{ 1,2,3 } , \
 '{ 1,2,7 } , \
 '{ 5,6,7 } , \
 '{ 2,3,7 } , \
 '{ 3,5,6 } , \
 '{ 1,2,7 } , \
 '{ 3,6,7 } , \
 '{ 1,2,3 } , \
 '{ 3,5,7 } , \
 '{ 1,2,3 } , \
 '{ 2,6,7 } , \
 '{ 1,3,6 } , \
 '{ 5,6,7 } , \
 '{ 1,6,7 } , \
 '{ 5,6,7 } , \
 '{ 5,6,7 } , \
 '{ 3,5,7 } , \
 '{ 2,3,6 } , \
 '{ 1,2,3 } , \
 '{ 2,3,5 } , \
 '{ 5,6,7 } , \
 '{ 3,5,7 } , \
 '{ 5,6,7 } , \
 '{ 2,5,7 } , \
 '{ 5,6,7 } , \
 '{ 3,5,6 } , \
 '{ 1,2,3 } , \
 '{ 1,2,3 } , \
 '{ 2,5,7 } , \
 '{ 1,3,6 }  }

`define TRIPLET_ADDER_DELAYS '{ \
 '{ 4,7,4 } , \
 '{ 21,23,27 } , \
 '{ 32,32,40 } , \
 '{ 17,18,19 } , \
 '{ 9,8,7 } , \
 '{ 17,17,15 } , \
 '{ 23,26,29 } , \
 '{ 18,19,20 } , \
 '{ 15,16,15 } , \
 '{ 29,28,32 } , \
 '{ 25,29,32 } , \
 '{ 31,35,28 } , \
 '{ 14,15,15 } , \
 '{ 27,32,36 } , \
 '{ 16,15,16 } , \
 '{ 34,44,39 } , \
 '{ 23,25,25 } , \
 '{ 11,10,10 } , \
 '{ 5,3,1 } , \
 '{ 19,21,23 } , \
 '{ 25,28,31 } , \
 '{ 34,34,38 } , \
 '{ 5,3,1 } , \
 '{ 9,8,7 } , \
 '{ 4,2,0 } , \
 '{ 17,18,19 } , \
 '{ 27,31,34 } , \
 '{ 20,22,24 } , \
 '{ 32,37,37 } , \
 '{ 15,15,14 } , \
 '{ 10,11,10 } , \
 '{ 26,30,33 } , \
 '{ 16,18,18 } , \
 '{ 26,22,24 } , \
 '{ 5,6,3 } , \
 '{ 8,7,6 } , \
 '{ 30,38,30 } , \
 '{ 19,21,23 } , \
 '{ 22,24,26 } , \
 '{ 18,19,20 } , \
 '{ 33,37,36 } , \
 '{ 27,21,23 } , \
 '{ 13,14,15 } , \
 '{ 16,16,16 } , \
 '{ 9,9,8 } , \
 '{ 41,32,41 } , \
 '{ 4,2,0 } , \
 '{ 34,35,39 } , \
 '{ 7,4,4 } , \
 '{ 21,23,25 } , \
 '{ 28,31,35 } , \
 '{ 25,28,31 } , \
 '{ 13,13,13 } , \
 '{ 42,32,42 } , \
 '{ 37,41,36 } , \
 '{ 11,11,11 } , \
 '{ 16,17,17 } , \
 '{ 12,12,12 } , \
 '{ 28,23,28 } , \
 '{ 10,10,9 } , \
 '{ 11,10,9 } , \
 '{ 24,27,30 } , \
 '{ 15,13,14 } , \
 '{ 13,13,13 } , \
 '{ 8,7,6 } , \
 '{ 39,34,44 } , \
 '{ 6,3,5 }  }

`define DOUBLET_ADDER_INDICES '{ \
 '{ 0,4  } , \
 '{ 0,4  } , \
 '{ 0,4  } , \
 '{ 0,4  } , \
 '{ 0,4  } , \
 '{ 0,4  } , \
 '{ 0,4  } , \
 '{ 0,4  } , \
 '{ 0,4  } , \
 '{ 0,4  } , \
 '{ 0,4  } , \
 '{ 0,4  }  }

`define DOUBLET_ADDER_DELAYS '{ \
 '{ 2,0  } , \
 '{ 1,0  } , \
 '{ 0,0  } , \
 '{ 4,1  } , \
 '{ 2,0  } , \
 '{ 4,0  } , \
 '{ 0,1  } , \
 '{ 2,1  } , \
 '{ 5,1  } , \
 '{ 3,0  } , \
 '{ 3,0  } , \
 '{ 1,1  }  }

`define BEAM_CONTENTS '{ \
 '{ 46,24,3 } , \
 '{ 34,66,3 } , \
 '{ 64,35,3 } , \
 '{ 23,4,1 } , \
 '{ 30,17,1 } , \
 '{ 63,52,1 } , \
 '{ 43,8,11 } , \
 '{ 25,3,11 } , \
 '{ 37,19,11 } , \
 '{ 38,33,11 } , \
 '{ 58,16,6 } , \
 '{ 51,20,6 } , \
 '{ 50,11,10 } , \
 '{ 21,36,10 } , \
 '{ 45,28,5 } , \
 '{ 65,15,5 } , \
 '{ 46,22,9 } , \
 '{ 66,0,9 } , \
 '{ 4,64,9 } , \
 '{ 44,59,0 } , \
 '{ 55,57,0 } , \
 '{ 42,12,0 } , \
 '{ 56,32,11 } , \
 '{ 39,3,2 } , \
 '{ 49,27,11 } , \
 '{ 1,33,6 } , \
 '{ 6,61,6 } , \
 '{ 10,31,6 } , \
 '{ 13,11,4 } , \
 '{ 36,47,4 } , \
 '{ 53,28,10 } , \
 '{ 18,24,9 } , \
 '{ 48,34,7 } , \
 '{ 23,35,7 } , \
 '{ 17,60,7 } , \
 '{ 63,57,7 } , \
 '{ 62,29,11 } , \
 '{ 5,14,2 } , \
 '{ 25,7,2 } , \
 '{ 27,19,6 } , \
 '{ 38,41,6 } , \
 '{ 61,20,4 } , \
 '{ 26,31,10 } , \
 '{ 9,40,10 } , \
 '{ 2,54,8 } , \
 '{ 65,15,8 }  }

