`define USING_DEBUG 0