`define BEAM_ANTENNA_DELAYS '{ \
	'{1,4,2,0,4,4,2,0}, \ // Beam 0
	'{0,5,4,2,3,5,4,2}, \ // Beam 1
	'{0,7,6,5,3,7,6,5}, \ // Beam 2
	'{0,9,8,7,1,9,8,7}, \ // Beam 3
	'{0,11,10,10,1,11,10,10}, \ // Beam 4
	'{0,13,13,13,1,13,13,13}, \ // Beam 5
	'{0,14,15,15,0,14,15,15}, \ // Beam 6
	'{0,16,17,18,0,16,17,18}, \ // Beam 7
	'{0,18,20,22,0,18,20,22}, \ // Beam 8
	'{0,21,23,25,0,21,23,25}, \ // Beam 9
	'{1,23,25,28,0,23,25,28}, \ // Beam 10
	'{1,25,28,31,0,25,28,31}, \ // Beam 11
	'{3,28,31,35,0,28,31,35}, \ // Beam 12
	'{3,30,34,38,0,30,34,38}, \ // Beam 13
	'{4,32,37,41,0,32,37,41}, \ // Beam 14
	'{4,34,39,44,0,34,39,44}, \ // Beam 15
	'{0,4,2,0,3,5,3,1}, \ // Beam 16
	'{0,6,4,3,3,7,5,4}, \ // Beam 17
	'{0,8,7,6,3,9,8,7}, \ // Beam 18
	'{0,9,9,8,2,10,10,9}, \ // Beam 19
	'{0,11,11,11,2,12,12,12}, \ // Beam 20
	'{0,13,14,14,2,15,15,15}, \ // Beam 21
	'{0,15,15,16,0,16,17,17}, \ // Beam 22
	'{0,17,18,19,0,18,19,20}, \ // Beam 23
	'{0,19,21,23,0,20,22,24}, \ // Beam 24
	'{1,21,23,26,0,22,24,27}, \ // Beam 25
	'{1,23,26,29,0,24,27,30}, \ // Beam 26
	'{1,25,29,32,0,26,30,33}, \ // Beam 27
	'{2,27,31,35,0,28,32,36}, \ // Beam 28
	'{2,30,34,38,0,30,35,39}, \ // Beam 29
	'{3,32,37,42,0,32,37,42}, \ // Beam 30
	'{0,5,3,1,3,4,2,0}, \ // Beam 31
	'{0,6,4,3,1,5,3,2}, \ // Beam 32
	'{0,8,7,6,1,7,6,5}, \ // Beam 33
	'{0,10,10,9,1,9,9,8}, \ // Beam 34
	'{0,12,12,12,1,11,11,11}, \ // Beam 35
	'{0,14,14,14,0,12,13,13}, \ // Beam 36
	'{0,16,17,17,0,15,15,16}, \ // Beam 37
	'{0,18,19,20,0,17,18,19}, \ // Beam 38
	'{1,20,22,24,0,19,21,23}, \ // Beam 39
	'{1,22,24,27,0,21,23,26}, \ // Beam 40
	'{2,25,28,31,0,24,27,30}, \ // Beam 41
	'{3,27,31,34,0,26,30,33}, \ // Beam 42
	'{3,29,33,37,0,28,32,36}, \ // Beam 43
	'{4,31,36,40,0,31,35,39}, \ // Beam 44
	'{4,33,38,43,0,33,38,43} \ // Beam 46
}
`define BEAM_TOTAL 46
`define MAX_ANTENNA_DELAY_0 4
`define MAX_ANTENNA_DELAY_1 34
`define MAX_ANTENNA_DELAY_2 39
`define MAX_ANTENNA_DELAY_3 44
`define MAX_ANTENNA_DELAY_4 4
`define MAX_ANTENNA_DELAY_5 34
`define MAX_ANTENNA_DELAY_6 39
`define MAX_ANTENNA_DELAY_7 44
