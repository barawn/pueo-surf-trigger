//`define BEAM_ANTENNA_DELAYS '{ '{1,4,2,0,4,4,2,0}, '{0,5,4,2,3,5,4,2}, '{0,7,6,5,3,7,6,5}, '{0,9,8,7,1,9,8,7}, '{0,11,10,10,1,11,10,10}, '{0,13,13,13,1,13,13,13}, '{0,14,15,15,0,14,15,15}, '{0,16,17,18,0,16,17,18}, '{0,18,20,22,0,18,20,22}, '{0,21,23,25,0,21,23,25}, '{1,23,25,28,0,23,25,28}, '{1,25,28,31,0,25,28,31}, '{3,28,31,35,0,28,31,35}, '{3,30,34,38,0,30,34,38}, '{4,32,37,41,0,32,37,41}, '{4,34,39,44,0,34,39,44}, '{0,4,2,0,3,5,3,1}, '{0,6,4,3,3,7,5,4}, '{0,8,7,6,3,9,8,7}, '{0,9,9,8,2,10,10,9}, '{0,11,11,11,2,12,12,12}, '{0,13,14,14,2,15,15,15}, '{0,15,15,16,0,16,17,17}, '{0,17,18,19,0,18,19,20}, '{0,19,21,23,0,20,22,24}, '{1,21,23,26,0,22,24,27}, '{1,23,26,29,0,24,27,30}, '{1,25,29,32,0,26,30,33}, '{2,27,31,35,0,28,32,36}, '{2,30,34,38,0,30,35,39}, '{3,32,37,42,0,32,37,42}, '{0,5,3,1,3,4,2,0}, '{0,6,4,3,1,5,3,2}, '{0,8,7,6,1,7,6,5}, '{0,10,10,9,1,9,9,8}, '{0,12,12,12,1,11,11,11}, '{0,14,14,14,0,12,13,13}, '{0,16,17,17,0,15,15,16}, '{0,18,19,20,0,17,18,19}, '{1,20,22,24,0,19,21,23}, '{1,22,24,27,0,21,23,26}, '{2,25,28,31,0,24,27,30}, '{3,27,31,34,0,26,30,33}, '{3,29,33,37,0,28,32,36}, '{4,31,36,40,0,31,35,39}, '{4,33,38,43,0,33,38,43} }
//`define FAKE_ANTENNA_DELAYS '{ '{0,0,0,0,0,0,0,0}, '{0,5,4,2,3,5,4,2}, '{0,7,6,5,3,7,6,5}, '{0,9,8,7,1,9,8,7}, '{0,11,10,10,1,11,10,10}, '{0,13,13,13,1,13,13,13}, '{0,14,15,15,0,14,15,15}, '{0,16,17,18,0,16,17,18}, '{0,18,20,22,0,18,20,22}, '{0,21,23,25,0,21,23,25}, '{1,23,25,28,0,23,25,28}, '{1,25,28,31,0,25,28,31}, '{3,28,31,35,0,28,31,35}, '{3,30,34,38,0,30,34,38}, '{4,32,37,41,0,32,37,41}, '{4,34,39,44,0,34,39,44}, '{0,4,2,0,3,5,3,1}, '{0,6,4,3,3,7,5,4}, '{0,8,7,6,3,9,8,7}, '{0,9,9,8,2,10,10,9}, '{0,11,11,11,2,12,12,12}, '{0,13,14,14,2,15,15,15}, '{0,15,15,16,0,16,17,17}, '{0,17,18,19,0,18,19,20}, '{0,19,21,23,0,20,22,24}, '{1,21,23,26,0,22,24,27}, '{1,23,26,29,0,24,27,30}, '{1,25,29,32,0,26,30,33}, '{2,27,31,35,0,28,32,36}, '{2,30,34,38,0,30,35,39}, '{3,32,37,42,0,32,37,42}, '{0,5,3,1,3,4,2,0}, '{0,6,4,3,1,5,3,2}, '{0,8,7,6,1,7,6,5}, '{0,10,10,9,1,9,9,8}, '{0,12,12,12,1,11,11,11}, '{0,14,14,14,0,12,13,13}, '{0,16,17,17,0,15,15,16}, '{0,18,19,20,0,17,18,19}, '{1,20,22,24,0,19,21,23}, '{1,22,24,27,0,21,23,26}, '{2,25,28,31,0,24,27,30}, '{3,27,31,34,0,26,30,33}, '{3,29,33,37,0,28,32,36}, '{4,31,36,40,0,31,35,39}, '{4,33,38,43,0,33,38,43} }
//`define BEAM_TOTAL 46
//`define MAX_ANTENNA_DELAY_0 4
//`define MAX_ANTENNA_DELAY_1 34
//`define MAX_ANTENNA_DELAY_2 39
//`define MAX_ANTENNA_DELAY_3 44
//`define MAX_ANTENNA_DELAY_4 4
//`define MAX_ANTENNA_DELAY_5 34
//`define MAX_ANTENNA_DELAY_6 39
//`define MAX_ANTENNA_DELAY_7 44

`define BEAM_ANTENNA_DELAYS '{'{4,0,-14,0,-36,-46,0,0},     \
                              '{1,0,-15,0,-38,-48,0,0},     \
                              '{0,1,-13,0,-10,-20,0,0},     \
                              '{4,0,-12,0,-33,-41,0,0},     \
                              '{1,0,-13,0,-35,-43,0,0},     \
                              '{0,1,-11,0,-7,-16,0,0},      \
                              '{4,0,-11,0,-29,-36,0,0},     \
                              '{0,0,-11,0,-31,-38,0,0},     \
                              '{0,0,-11,0,-6,-13,0,0},      \
                              '{0,1,-13,0,-36,0,-48,0}, '{0,4,-10,0,-32,0,-46,0}, '{1,0,-15,0,-11,0,-20,0}, '{4,0,-14,0,-13,0,-19,0}, '{0,1,-11,0,-33,0,-43,0}, '{0,4,-9,0,-29,0,-41,0}, '{1,0,-13,0,-9,0,-16,0}, '{4,0,-12,0,-10,0,-15,0}, '{0,4,-8,0,-26,0,-36,0}, '{4,0,-11,0,-7,0,-11,0}, '{0,0,-14,-16,0,0,-49,-48}, '{0,0,-14,-13,0,0,-47,-48}, '{0,0,-14,-10,0,0,-42,-46}, '{0,0,-14,-13,0,0,-20,-21}, '{0,0,-14,-16,0,0,-23,-21}, '{0,0,-13,-14,0,0,-44,-43}, '{0,0,-13,-11,0,0,-42,-43}, '{0,0,-13,-9,0,0,-38,-41}, '{0,0,-13,-11,0,0,-16,-17}, '{0,0,-13,-14,0,0,-18,-17}, '{0,0,-11,-11,0,0,-38,-38}, '{0,0,-11,-8,0,0,-33,-36}, '{0,0,-11,-11,0,0,-13,-13}, '{0,0,0,-1,-12,-23,0,-36}, '{0,0,0,-1,-10,-20,0,-33}, '{0,0,0,-2,-9,-19,0,-31}, '{0,0,0,-26,-32,-42,0,-31}, '{0,0,0,-28,-36,-47,0,-33}, '{0,0,0,-28,-39,-49,0,-36}, '{0,0,0,0,-10,-18,0,-31}, '{0,0,0,0,-7,-16,0,-29}, '{0,0,0,-1,-6,-15,0,-26}, '{0,0,0,-24,-29,-38,0,-26}, '{0,0,0,-26,-33,-42,0,-29}, '{0,0,0,-26,-36,-44,0,-31}, '{0,0,0,1,-6,-13,0,-26}, '{0,0,0,-1,-4,-11,0,-22}, '{0,0,0,-22,-26,-33,0,-22}, '{0,0,0,-24,-31,-38,0,-26} }

`define BEAM_USED_CHANNELS '{8'b11101100,       \
                             8'b11101100,       \
                             8'b11101100,       \
                             8'b11101100,       \
                             8'b11101100,       \
                             8'b11101100,       \
                             8'b11101100,       \
                             8'b11101100,       \
                             8'b11101100,       \
                             8'b11101010, 8'b11101010, 8'b11101010, 8'b11101010, 8'b11101010, 8'b11101010, 8'b11101010, 8'b11101010, 8'b11101010, 8'b11101010, 8'b01110011, 8'b01110011, 8'b01110011, 8'b01110011, 8'b01110011, 8'b01110011, 8'b01110011, 8'b01110011, 8'b01110011, 8'b01110011, 8'b01110011, 8'b01110011, 8'b01110011, 8'b10011101, 8'b10011101, 8'b10011101, 8'b10011101, 8'b10011101, 8'b10011101, 8'b10011101, 8'b10011101, 8'b10011101, 8'b10011101, 8'b10011101, 8'b10011101, 8'b10011101, 8'b10011101, 8'b10011101, 8'b10011101}

`define BEAM_CHANNEL_INVERSION '{8'b00001100,   \
                                 8'b00001100,   \
                                 8'b11100000,   \
                                 8'b00001100,   \
                                 8'b00001100,   \
                                 8'b11100000,   \
                                 8'b00001100,   \
                                 8'b00001100,   \
                                 8'b11100000,   \
                                 8'b00001010, 8'b00001010, 8'b11100000, 8'b11100000, 8'b00001010, 8'b00001010, 8'b11100000, 8'b11100000, 8'b00001010, 8'b11100000, 8'b00000011, 8'b00000011, 8'b00000011, 8'b01110000, 8'b01110000, 8'b00000011, 8'b00000011, 8'b00000011, 8'b01110000, 8'b01110000, 8'b00000011, 8'b00000011, 8'b01110000, 8'b10000001, 8'b10000001, 8'b10000001, 8'b00011100, 8'b00011100, 8'b00011100, 8'b10000001, 8'b10000001, 8'b10000001, 8'b00011100, 8'b00011100, 8'b00011100, 8'b10000001, 8'b10000001, 8'b00011100, 8'b00011100 }

//for TEB0835 testing we only have access to 0,2,4,6
//`define BEAM_ANTENNA_DELAYS '{'{4,0,0,0,-16,0,-39,-51}, '{1,0,-16,0,-41,-53,0,0}}
//`define BEAM_ANTENNA_DELAYS '{'{0,0,4,0,20,0,43,55}, '{1,0,-16,0,-41,-53,0,0}}
//`define BEAM_ANTENNA_DELAYS '{'{0,0,0,0,0,0,0,0}, '{1,0,-16,0,-41,-53,0,0}}
//`define BEAM_USED_CHANNELS '{8'b10101011, 8'b11101100}
//`define BEAM_CHANNEL_INVERSION '{8'b00000011, 8'b00001100}

`define BEAM_TOTAL 48
`define MAX_ANTENNA_DELAY_0 4
`define MAX_ANTENNA_DELAY_1 34
`define MAX_ANTENNA_DELAY_2 39
`define MAX_ANTENNA_DELAY_3 44
`define MAX_ANTENNA_DELAY_4 4
`define MAX_ANTENNA_DELAY_5 34
`define MAX_ANTENNA_DELAY_6 39
`define MAX_ANTENNA_DELAY_7 44
