`ifndef PUEO_LF_META_SV
`define PUEO_LF_META_SV

package pueo_lf_meta;

   localparam int LF_META7_INDICES [0:21] = ' {
	36,
	37,
	42,
	43,
	46,
	47,
	255,
	255,

	255,
	255,
	255,
	255,
	255,
	255,
	255,
	255,

	255,
	255,
	255,
	255,
	255,
	255};

   localparam int LF_META6_INDICES [0:21] = ' {
	23,
	27,
	28,
	31,
	35,
	41,
	255,
	255,

	255,
	255,
	255,
	255,
	255,
	255,
	255,
	255,

	255,
	255,
	255,
	255,
	255,
	255 };


   localparam int LF_META5_INDICES [0:21] = ' {
	11,
	12,
	15,
	16,
	18,
	22,
	255,
	255,

	255,
	255,
	255,
	255,
	255,
	255,
	255,
	255,

	255,
	255,
	255,
	255,
	255,
	255 };


   localparam int LF_META4_INDICES [0:21] = ' {
	2,
	5,
	8,
	34,
	40,
	45,
	255,
	255,

	255,
	255,
	255,
	255,
	255,
	255,
	255,
	255,

	255,
	255,
	255,
	255,
	255,
	255 };

   localparam int LF_META3_INDICES [0:21] = ' {
	30,
	32,
	33,
	38,
	39,
	44,
	255,
	255,

	255,
	255,
	255,
	255,
	255,
	255,
	255,
	255,

	255,
	255,
	255,
	255,
	255,
	255 };


   localparam int LF_META2_INDICES [0:21] = ' {
	20,
	21,
	24,
	25,
	26,
	29,
	255,
	255,

	255,
	255,
	255,
	255,
	255,
	255,
	255,
	255,

	255,
	255,
	255,
	255,
	255,
	255 };


   localparam int LF_META1_INDICES [0:21] = ' {
	9,
	10,
	13,
	14,
	17,
	19,
	255,
	255,

	255,
	255,
	255,
	255,
	255,
	255,
	255,
	255,

	255,
	255,
	255,
	255,
	255,
	255 };

   localparam int LF_META0_INDICES [0:21] = ' {
	0,
	1,
	3,
	4,
	6,
	7,
	255,
	255,

	255,
	255,
	255,
	255,
	255,
	255,
	255,
	255,

	255,
	255,
	255,
	255,
	255,
	255 };

endpackage // pueo_lf_meta

`endif
