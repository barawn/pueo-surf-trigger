//True beams
`define BEAM_ANTENNA_DELAYS '{'{-36,-46,0,0,4,0,-14,0}, '{-38,-48,0,0,1,0,-15,0}, '{-10,-20,0,0,0,1,-13,0}, '{-33,-41,0,0,4,0,-12,0}, '{-35,-43,0,0,1,0,-13,0}, '{-7,-16,0,0,0,1,-11,0}, '{-29,-36,0,0,4,0,-11,0}, '{-31,-38,0,0,0,0,-11,0}, '{-6,-13,0,0,0,0,-11,0}, '{-36,0,-48,0,0,1,-13,0}, '{-32,0,-46,0,0,4,-10,0}, '{-11,0,-20,0,1,0,-15,0}, '{-13,0,-19,0,4,0,-14,0}, '{-33,0,-43,0,0,1,-11,0}, '{-29,0,-41,0,0,4,-9,0}, '{-9,0,-16,0,1,0,-13,0}, '{-10,0,-15,0,4,0,-12,0}, '{-26,0,-36,0,0,4,-8,0}, '{-7,0,-11,0,4,0,-11,0}, '{0,0,-49,-48,0,0,-14,-16}, '{0,0,-47,-48,0,0,-14,-13}, '{0,0,-42,-46,0,0,-14,-10}, '{0,0,-20,-21,0,0,-14,-13}, '{0,0,-23,-21,0,0,-14,-16}, '{0,0,-44,-43,0,0,-13,-14}, '{0,0,-42,-43,0,0,-13,-11}, '{0,0,-38,-41,0,0,-13,-9}, '{0,0,-16,-17,0,0,-13,-11}, '{0,0,-18,-17,0,0,-13,-14}, '{0,0,-38,-38,0,0,-11,-11}, '{0,0,-33,-36,0,0,-11,-8}, '{0,0,-13,-13,0,0,-11,-11}, '{-12,-23,0,-36,0,0,0,-1}, '{-10,-20,0,-33,0,0,0,-1}, '{-9,-19,0,-31,0,0,0,-2}, '{-32,-42,0,-31,0,0,0,-26}, '{-36,-47,0,-33,0,0,0,-28}, '{-39,-49,0,-36,0,0,0,-28}, '{-10,-18,0,-31,0,0,0,0}, '{-7,-16,0,-29,0,0,0,0}, '{-6,-15,0,-26,0,0,0,-1}, '{-29,-38,0,-26,0,0,0,-24}, '{-33,-42,0,-29,0,0,0,-26}, '{-36,-44,0,-31,0,0,0,-26}, '{-6,-13,0,-26,0,0,0,1}, '{-4,-11,0,-22,0,0,0,-1}, '{-26,-33,0,-22,0,0,0,-22}, '{-31,-38,0,-26,0,0,0,-24} }
`define BEAM_USED_CHANNELS '{8'b11001110, 8'b11001110, 8'b11001110, 8'b11001110, 8'b11001110, 8'b11001110, 8'b11001110, 8'b11001110, 8'b11001110, 8'b10101110, 8'b10101110, 8'b10101110, 8'b10101110, 8'b10101110, 8'b10101110, 8'b10101110, 8'b10101110, 8'b10101110, 8'b10101110, 8'b00110111, 8'b00110111, 8'b00110111, 8'b00110111, 8'b00110111, 8'b00110111, 8'b00110111, 8'b00110111, 8'b00110111, 8'b00110111, 8'b00110111, 8'b00110111, 8'b00110111, 8'b11011001, 8'b11011001, 8'b11011001, 8'b11011001, 8'b11011001, 8'b11011001, 8'b11011001, 8'b11011001, 8'b11011001, 8'b11011001, 8'b11011001, 8'b11011001, 8'b11011001, 8'b11011001, 8'b11011001, 8'b11011001}
//For HPOLE compile
`define BEAM_CHANNEL_INVERSION '{8'b11000000, 8'b11000000, 8'b00001110, 8'b11000000, 8'b11000000, 8'b00001110, 8'b11000000, 8'b11000000, 8'b00001110, 8'b10100000, 8'b10100000, 8'b00001110, 8'b00001110, 8'b10100000, 8'b10100000, 8'b00001110, 8'b00001110, 8'b10100000, 8'b00001110, 8'b00110000, 8'b00110000, 8'b00110000, 8'b00000111, 8'b00000111, 8'b00110000, 8'b00110000, 8'b00110000, 8'b00000111, 8'b00000111, 8'b00110000, 8'b00110000, 8'b00000111, 8'b00011000, 8'b00011000, 8'b00011000, 8'b11000001, 8'b11000001, 8'b11000001, 8'b00011000, 8'b00011000, 8'b00011000, 8'b11000001, 8'b11000001, 8'b11000001, 8'b00011000, 8'b00011000, 8'b11000001, 8'b11000001}
//For VPOLE compile
//`define BEAM_CHANNEL_INVERSION '{8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000}

//new beamforming - not in use
//`define BEAM_ANTENNA_DELAYS '{'{-36,-46,0,0,4,0,-14,0}, '{-38,-48,0,0,1,0,-15,0}, '{-10,-20,0,0,0,1,-13,0}, '{-33,-41,0,0,4,0,-12,0}, '{-35,-43,0,0,1,0,-13,0}, '{-7,-16,0,0,0,1,-11,0}, '{-29,-36,0,0,4,0,-11,0}, '{-31,-38,0,0,0,0,-11,0}, '{-6,-13,0,0,0,0,-11,0}, '{-36,0,-48,0,0,1,-13,0}, '{-32,0,-46,0,0,4,-10,0}, '{-11,0,-20,0,1,0,-15,0}, '{-13,0,-19,0,4,0,-14,0}, '{-33,0,-43,0,0,1,-11,0}, '{-29,0,-41,0,0,4,-9,0}, '{-9,0,-16,0,1,0,-13,0}, '{-10,0,-15,0,4,0,-12,0}, '{-26,0,-36,0,0,4,-8,0}, '{-7,0,-11,0,4,0,-11,0}, '{0,0,-49,-48,0,0,-14,-16}, '{0,0,-47,-48,0,0,-14,-13}, '{0,0,-42,-46,0,0,-14,-10}, '{0,0,-20,-21,0,0,-14,-13}, '{0,0,-23,-21,0,0,-14,-16}, '{0,0,-44,-43,0,0,-13,-14}, '{0,0,-42,-43,0,0,-13,-11}, '{0,0,-38,-41,0,0,-13,-9}, '{0,0,-16,-17,0,0,-13,-11}, '{0,0,-18,-17,0,0,-13,-14}, '{0,0,-38,-38,0,0,-11,-11}, '{0,0,-33,-36,0,0,-11,-8}, '{0,0,-13,-13,0,0,-11,-11}, '{-12,-23,0,-36,0,0,0,-1}, '{-10,-20,0,-33,0,0,0,-1}, '{-9,-19,0,-31,0,0,0,-2}, '{-32,-42,0,-31,0,0,0,-26}, '{-36,-47,0,-33,0,0,0,-28}, '{-39,-49,0,-36,0,0,0,-28}, '{-10,-18,0,-31,0,0,0,0}, '{-7,-16,0,-29,0,0,0,0}, '{-6,-15,0,-26,0,0,0,-1}, '{-29,-38,0,-26,0,0,0,-24}, '{-33,-42,0,-29,0,0,0,-26}, '{-36,-44,0,-31,0,0,0,-26}, '{-6,-13,0,-26,0,0,0,1}, '{-4,-11,0,-22,0,0,0,-1}, '{-26,-33,0,-22,0,0,0,-22}, '{-31,-38,0,-26,0,0,0,-24} }
//`define BEAM_USED_CHANNELS '{ '{0,1,4,5,6},  '{0,1,4,5,6},  '{0,1,4,5,6},  '{0,1,4,5,6},  '{0,1,4,5,6},  '{0,1,4,5,6},  '{0,1,4,5,6},  '{0,1,4,5,6},  '{0,1,4,5,6},  '{0,2,4,5,6},  '{0,2,4,5,6},  '{0,2,4,5,6},  '{0,2,4,5,6},  '{0,2,4,5,6},  '{0,2,4,5,6},  '{0,2,4,5,6},  '{0,2,4,5,6},  '{0,2,4,5,6},  '{0,2,4,5,6},  '{2,3,5,6,7},  '{2,3,5,6,7},  '{2,3,5,6,7},  '{2,3,5,6,7},  '{2,3,5,6,7},  '{2,3,5,6,7},  '{2,3,5,6,7},  '{2,3,5,6,7},  '{2,3,5,6,7},  '{2,3,5,6,7},  '{2,3,5,6,7},  '{2,3,5,6,7},  '{2,3,5,6,7},  '{0,1,3,4,7},  '{0,1,3,4,7},  '{0,1,3,4,7},  '{0,1,3,4,7},  '{0,1,3,4,7},  '{0,1,3,4,7},  '{0,1,3,4,7},  '{0,1,3,4,7},  '{0,1,3,4,7},  '{0,1,3,4,7},  '{0,1,3,4,7},  '{0,1,3,4,7},  '{0,1,3,4,7},  '{0,1,3,4,7},  '{0,1,3,4,7},  '{0,1,3,4,7}}
//For HPOLE compile
//`define BEAM_CHANNEL_INVERSION '{ '{1,1,0,0,0}, '{1,1,0,0,0}, '{0,0,1,1,1}, '{1,1,0,0,0}, '{1,1,0,0,0}, '{0,0,1,1,1}, '{1,1,0,0,0}, '{1,1,0,0,0}, '{0,0,1,1,1}, '{1,1,0,0,0}, '{1,1,0,0,0}, '{0,0,1,1,1}, '{0,0,1,1,1}, '{1,1,0,0,0}, '{1,1,0,0,0}, '{0,0,1,1,1}, '{0,0,1,1,1}, '{1,1,0,0,0}, '{0,0,1,1,1}, '{1,1,0,0,0}, '{1,1,0,0,0}, '{1,1,0,0,0}, '{0,0,1,1,1}, '{0,0,1,1,1}, '{1,1,0,0,0}, '{1,1,0,0,0}, '{1,1,0,0,0}, '{0,0,1,1,1}, '{0,0,1,1,1}, '{1,1,0,0,0}, '{1,1,0,0,0}, '{0,0,1,1,1}, '{0,0,1,1,0}, '{0,0,1,1,0}, '{0,0,1,1,0}, '{1,1,0,0,1}, '{1,1,0,0,1}, '{1,1,0,0,1}, '{0,0,1,1,0}, '{0,0,1,1,0}, '{0,0,1,1,0}, '{1,1,0,0,1}, '{1,1,0,0,1}, '{1,1,0,0,1}, '{0,0,1,1,0}, '{0,0,1,1,0}, '{1,1,0,0,1}, '{1,1,0,0,1}}
//For VPOLE compile
//`define BEAM_CHANNEL_INVERSION '{ '{0,0,0,0,0}, '{0,0,0,0,0}, '{0,0,0,0,0}, '{0,0,0,0,0}, '{0,0,0,0,0}, '{0,0,0,0,0}, '{0,0,0,0,0}, '{0,0,0,0,0}, '{0,0,0,0,0}, '{0,0,0,0,0}, '{0,0,0,0,0}, '{0,0,0,0,0}, '{0,0,0,0,0}, '{0,0,0,0,0}, '{0,0,0,0,0}, '{0,0,0,0,0}, '{0,0,0,0,0}, '{0,0,0,0,0}, '{0,0,0,0,0}, '{0,0,0,0,0}, '{0,0,0,0,0}, '{0,0,0,0,0}, '{0,0,0,0,0}, '{0,0,0,0,0}, '{0,0,0,0,0}, '{0,0,0,0,0}, '{0,0,0,0,0}, '{0,0,0,0,0}, '{0,0,0,0,0}, '{0,0,0,0,0}, '{0,0,0,0,0}, '{0,0,0,0,0}, '{0,0,0,0,0}, '{0,0,0,0,0}, '{0,0,0,0,0}, '{0,0,0,0,0}, '{0,0,0,0,0}, '{0,0,0,0,0}, '{0,0,0,0,0}, '{0,0,0,0,0}, '{0,0,0,0,0}, '{0,0,0,0,0}, '{0,0,0,0,0}, '{0,0,0,0,0}, '{0,0,0,0,0}, '{0,0,0,0,0}, '{0,0,0,0,0}, '{0,0,0,0,0}}


//for TEB0835 testing we only have access to 0,2,4,6
//`define BEAM_ANTENNA_DELAYS '{'{4,0,0,0,-14,0,-36,0}, '{1,0,0,0,-15,0,-38,0}, '{0,0,1,0,-13,0,-10,0}, '{4,0,0,0,-12,0,-33,0}, '{1,0,0,0,-13,0,-35,0}, '{0,0,1,0,-11,0,-7,0}, '{4,0,0,0,-11,0,-29,0}, '{0,0,0,0,-11,0,-31,0}, '{0,0,0,0,-11,0,-6,0}, '{0,0,1,0,-13,0,-36,0}, '{0,0,4,0,-10,0,-32,0}, '{1,0,0,0,-15,0,-11,0}, '{4,0,0,0,-14,0,-13,0}, '{0,0,1,0,-11,0,-33,0}, '{0,0,4,0,-9,0,-29,0}, '{1,0,0,0,-13,0,-9,0}, '{4,0,0,0,-12,0,-10,0}, '{0,0,4,0,-8,0,-26,0}, '{4,0,0,0,-11,0,-7,0}, '{0,0,-14,0,-16,0,-49,0}, '{0,0,-14,0,-13,0,-47,0}, '{0,0,-14,0,-10,0,-42,0}, '{0,0,-14,0,-13,0,-20,0}, '{0,0,-14,0,-16,0,-23,0}, '{0,0,-13,0,-14,0,-44,0}, '{0,0,-13,0,-11,0,-42,0}, '{0,0,-13,0,-9,0,-38,0}, '{0,0,-13,0,-11,0,-16,0}, '{0,0,-13,0,-14,0,-18,0}, '{0,0,-11,0,-11,0,-38,0}, '{0,0,-11,0,-8,0,-33,0}, '{0,0,-11,0,-11,0,-13,0}, '{0,0,-1,0,-12,0,-23,0}, '{0,0,-1,0,-10,0,-20,0}, '{0,0,-2,0,-9,0,-19,0}, '{0,0,-26,0,-32,0,-42,0}, '{0,0,-28,0,-36,0,-47,0}, '{0,0,-28,0,-39,0,-49,0}, '{0,0,0,0,-10,0,-18,0}, '{0,0,0,0,-7,0,-16,0}, '{0,0,-1,0,-6,0,-15,0}, '{0,0,-24,0,-29,0,-38,0}, '{0,0,-26,0,-33,0,-42,0}, '{0,0,-26,0,-36,0,-44,0}, '{0,0,1,0,-6,0,-13,0}, '{0,0,-1,0,-4,0,-11,0}, '{0,0,-22,0,-26,0,-33,0}, '{0,0,-24,0,-31,0,-38,0}}
//`define BEAM_ANTENNA_DELAYS '{'{0,0,4,0,20,0,43,55}, '{1,0,-16,0,-41,-53,0,0}}
//`define BEAM_ANTENNA_DELAYS '{'{0,0,0,0,0,0,0,0}, '{1,0,-16,0,-41,-53,0,0}}
//OLD

//`define BEAM_USED_CHANNELS '{8'b10101011,8'b10101011,8'b10101011,8'b10101011,8'b10101011,8'b10101011,8'b10101011,8'b10101011,8'b10101011,8'b10101011,8'b10101011,8'b10101011,8'b10101011,8'b10101011,8'b10101011,8'b10101011,8'b10101011,8'b10101011,8'b10101011,8'b10101011,8'b10101011,8'b10101011,8'b10101011,8'b10101011,8'b10101011,8'b10101011,8'b10101011,8'b10101011,8'b10101011,8'b10101011,8'b10101011,8'b10101011,8'b10101011,8'b10101011,8'b10101011,8'b10101011,8'b10101011,8'b10101011,8'b10101011,8'b10101011,8'b10101011,8'b10101011,8'b10101011,8'b10101011,8'b10101011,8'b10101011,8'b10101011,8'b10101011}
//`define BEAM_CHANNEL_INVERSION '{8'b00000010, 8'b00000010, 8'b10101000, 8'b00000010, 8'b00000010, 8'b10101000, 8'b00000010, 8'b00000010, 8'b10101000, 8'b00000010, 8'b00000010, 8'b10101000, 8'b10101000, 8'b00000010, 8'b00000010, 8'b10101000, 8'b10101000, 8'b00000010, 8'b10101000, 8'b00000010, 8'b00000010, 8'b00000010, 8'b10101000, 8'b10101000, 8'b00000010, 8'b00000010, 8'b00000010, 8'b10101000, 8'b10101000, 8'b00000010, 8'b00000010, 8'b10101000, 8'b10000000, 8'b10000000, 8'b10000000, 8'b00101010, 8'b00101010, 8'b00101010, 8'b10000000, 8'b10000000, 8'b10000000, 8'b00101010, 8'b00101010, 8'b00101010, 8'b10000000, 8'b10000000, 8'b00101010, 8'b00101010}

`define BEAM_TOTAL 48
`define MAX_ANTENNA_DELAY_0 4
`define MAX_ANTENNA_DELAY_1 34
`define MAX_ANTENNA_DELAY_2 39
`define MAX_ANTENNA_DELAY_3 44
`define MAX_ANTENNA_DELAY_4 4
`define MAX_ANTENNA_DELAY_5 34
`define MAX_ANTENNA_DELAY_6 39
`define MAX_ANTENNA_DELAY_7 44
